class random_seq extends base_seq;


        `uvm_object_utils(ramdom_seq)

  //alu_config  m_config;

  extern function new(string name = "");
  extern task body();


endclass : base_seq


function base_seq::new(string name = "");
  super.new(name);
endfunction : new


task base_seq::body();
  `uvm_info(get_type_name(), "Random sequence starting", UVM_HIGH)
 
  repeat (5) begin

  req = apb_transaction::type_id::create("req");
  start_item(req); 
  if ( !req.randomize() )
    `uvm_error(get_type_name(), "Failed to randomize transaction")
  finish_item(req);
    
  end

  `uvm_info(get_type_name(), "Random sequence completed", UVM_HIGH)
endtask : body

`endif // BASE_SEQ_SV

