// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: top_test_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Fri Feb 13 17:50:22 2026
//=============================================================================
// Description: Test package for top
//=============================================================================

`ifndef TEST_PKG_SV
`define TEST_PKG_SV

package test_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;
  import env_pkg::*;

  `include "base_test.sv"

endpackage : test_pkg

`endif // TEST_PKG_SV

