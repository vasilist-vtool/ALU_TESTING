class driver extends uvm;

endclass
