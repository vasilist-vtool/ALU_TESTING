`ifndef ALU_SEQUENCER_SV
`define ALU_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(apb_transaction) alu_sequencer_t;


`endif // ALU_SEQUENCER_SV