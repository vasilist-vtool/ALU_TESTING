//Sequences
`include "sequences/base_seq.sv"