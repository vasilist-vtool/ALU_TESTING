package alu_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;
  import top_pkg::*;


`include "apb_transaction.sv"
`include "alu_config.sv"
`include "alu_driver.sv"
`include "alu_monitor.sv"
`include "alu_sequencer.sv"
//   `include "alu_coverage.sv"
`include "alu_agent.sv"
`include "alu_seq_lib.sv"

endpackage : alu_pkg
