

package env_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;

  `include "alu_env.sv"

endpackage : env_pkg

