//Sequences
`include "sequences/base_seq.sv"
`include "sequences/random_seq.sv"
`include "sequences/write_only_seq.sv"
`include "sequences/read_only_seq.sv"
