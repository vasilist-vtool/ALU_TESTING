
`ifndef ALU_IF_SV
`define ALU_IF_SV

interface alu_if(); 

  timeunit      1ns;
  timeprecision 1ps;

  //import alu_pkg::*;
  logic clk ;
  logic [`ADDR_W:0] paddr;
  logic [(`APB_BUS_SIZE-1):0] pwdata;
  logic [(`APB_BUS_SIZE-1):0] prdata;
  logic       penable;
  logic       pwrite;
  logic       psel;
  logic       rst_n;
  logic       ready;
  logic       slv_err;

  // You can insert properties and assertions here

endinterface : alu_if

`endif // ALU_IF_SV