package top_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;

  `include "defines.sv"


endpackage : top_pkg

