//Sequences
`include "sequences/base_seq.sv"
`include "sequences/random_seq.sv"