

package env_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;
  
  `include "virtual_sequence.sv"
  `include "alu_env.sv"

endpackage : env_pkg

