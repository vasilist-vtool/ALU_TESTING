`ifndef TEST_PKG_SV
`define TEST_PKG_SV

package test_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import alu_pkg::*;
  import env_pkg::*;

  `include "base_test.sv"

endpackage : test_pkg

`endif 

