`define DATA_WIDTH 16
`define DATA_SIZE 16
`define MUL_DATA_SIZE 8
`define FIFO_IN_DEPTH 4
`define FIFO_OUT_DEPTH 4
`define FIFO_IN_WIDTH 42
`define FIFO_OUT_WIDTH 25
`define APB_BUS_SIZE 32
`define REG_NUMBER 5
`define ADDR_W 2


typedef enum {read, write} wr_rd_type;

//for coverage
typedef enum {write_to_read_register,
              read_from_write_register,
              no_available_addr,
              read_from_empty_fifo_out,
              write_to_full_fifo_in,
              false_operation
} cause_of_slv_err;

typedef enum  { addition,
               multiplication
} operation_type;


typedef enum  { apb_write,
               apb_read_monitor,
               apb_read_slv_err,
               apb_read_no_slav_err,
               comparison_succesful
} checker_type;

typedef logic[`ADDR_W : 0] address_t;
typedef logic[`APB_BUS_SIZE-1 : 0] data_t;

typedef enum  { ALU_TX_STATE_IDLE,
                ALU_TX_STATE_ACTIVE,
                ALU_TX_STATE_COMPLETED
} alu_tx_state;

int NUM_TRANSACTIONS = 10;
int MAX_DELAY = 10;
int MIN_DELAY = 0;